module sega(W, X, Y, Z, OUT, OUTNAND);
  input  W;
  input  X;
  input  Y;
  input  Z;
  
  output OUT;
  output OUTNAND;
  

endmodule
